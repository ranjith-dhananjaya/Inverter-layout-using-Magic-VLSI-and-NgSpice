magic
tech scmos
timestamp 1640207986
<< nwell >>
rect -8 -1 10 17
<< polysilicon >>
rect 0 7 2 9
rect 0 -4 2 0
rect 1 -8 2 -4
rect 0 -11 2 -8
rect 0 -17 2 -15
<< ndiffusion >>
rect -2 -15 0 -11
rect 2 -15 3 -11
rect 7 -15 8 -11
<< pdiffusion >>
rect -6 5 0 7
rect -2 1 0 5
rect -6 0 0 1
rect 2 5 8 7
rect 2 1 3 5
rect 7 1 8 5
rect 2 0 8 1
<< metal1 >>
rect -2 12 3 16
rect 7 12 8 16
rect -5 5 -2 12
rect 4 5 7 6
rect 4 -4 7 1
rect -8 -8 -3 -4
rect 4 -8 14 -4
rect 4 -11 7 -8
rect -5 -20 -2 -15
rect -2 -24 3 -20
rect 7 -24 8 -20
<< ntransistor >>
rect 0 -15 2 -11
<< ptransistor >>
rect 0 0 2 7
<< polycontact >>
rect -3 -8 1 -4
<< ndcontact >>
rect -6 -15 -2 -11
rect 3 -15 7 -11
<< pdcontact >>
rect -6 1 -2 5
rect 3 1 7 5
<< psubstratepcontact >>
rect -6 -24 -2 -20
rect 3 -24 7 -20
<< nsubstratencontact >>
rect -6 12 -2 16
rect 3 12 7 16
<< labels >>
rlabel metal1 0 -22 0 -22 1 gnd
rlabel metal1 0 14 0 14 5 vdd
rlabel metal1 -8 -8 -8 -4 3 in
rlabel metal1 14 -8 14 -4 7 out
<< end >>
